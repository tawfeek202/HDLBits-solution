// todo A 32-bit vector can be viewed as containing 4 bytes (bits [31:24], [23:16], etc.). 
// todo Build a circuit that will reverse the byte ordering of the 4-byte word.
// todo AaaaaaaaBbbbbbbbCcccccccDddddddd => DdddddddCcccccccBbbbbbbbAaaaaaaa
module Vector2 (
    input  [31:0] in,
    output [31:0] out
);

  assign out[31 : 24] = in[7:0];
  assign out[23 : 16] = in[15:8];
  assign out[15 : 8]  = in[23:16];
  assign out[7 : 0]   = in[31:24];

endmodule

`timescale 1us / 1ns
module Wiredecl_TB ();

  /////////////////////////////////////////////////////////
  ///////////////////// Parameters ////////////////////////
  /////////////////////////////////////////////////////////

  parameter Clock_PERIOD = 10;

  /////////////////////////////////////////////////////////
  //////////////////// DUT Signals ////////////////////////
  /////////////////////////////////////////////////////////
  //*Inputs
  reg  a_TB;
  reg  b_TB;
  reg  c_TB;
  reg  d_TB;

  //* Outputs
  wire out_TB;
  wire out_n_TB;
  ////////////////////////////////////////////////////////
  ////////////////// initial block /////////////////////// 
  ////////////////////////////////////////////////////////


  initial begin
    //^ generating VCD file "value change dump"

    $dumpfile("Wiredecl.vcd");
    $dumpvars(0, Wiredecl_TB);

    ////////////////////////////////////////////////////////////////
    ///////////////////observing the wire output ///////////////////
    ////////////////////////////////////////////////////////////////

    //Note : out = (a & b) | (c & d) ;
    //Note : out_n = ~((a & b) | (c & d));

    //*apply all the scenarios you want




















  end
  ////////////////////////////////////////////////////////
  /////////////////// DUT Instantation ///////////////////
  ////////////////////////////////////////////////////////
  Wiredecl DUT (

      //*Inputs
      .a(a_TB),
      .b(b_TB),
      .c(c_TB),
      .d(d_TB),

      //* Outputs
      .out  (out_TB),
      .out_n(out_n_TB)
  );

endmodule

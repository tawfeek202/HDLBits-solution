`timescale 1us / 1ns
module ONE_TB ();

  /////////////////////////////////////////////////////////
  ///////////////////// Parameters ////////////////////////
  /////////////////////////////////////////////////////////

  parameter Clock_PERIOD = 10;

  /////////////////////////////////////////////////////////
  //////////////////// DUT Signals ////////////////////////
  /////////////////////////////////////////////////////////

  //* outputs
  wire one_TB;

  ////////////////////////////////////////////////////////
  ////////////////// initial block /////////////////////// 
  ////////////////////////////////////////////////////////


  initial begin
    //^ generating VCD file "value change dump"

    $dumpfile("ONE.vcd");
    $dumpvars(0, ONE_TB);

    ////////////////////////////////////////////////////////////////
    ///////////////////observing the output is one ///////////////////
    ////////////////////////////////////////////////////////////////

    $display("****************** one ***************");
    #Clock_PERIOD

      if (one_TB == 1) begin

        $display("test case succedded");

      end else begin

        $display("test case failed");

      end

  end
  ////////////////////////////////////////////////////////
  /////////////////// DUT Instantation ///////////////////
  ////////////////////////////////////////////////////////
  ONE DUT (
      //* Outputs
      .one(one_TB)
  );

endmodule

module ONE (
    output one
);
  assign one = 1'b1;
endmodule

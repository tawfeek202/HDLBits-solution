module NOT (
    input  in,
    output out
);
  assign out = ~in;
endmodule
